* MBR0520LT1G

.SUBCKT MBR0520LT1G A C
	* Connections
	D1 A C DMBR0520lT1

	.MODEL DMBR0520lT1 d
	+IS=1e-06 RS=0.115754 N=0.874519 EG=0.6
	+XTI=2.49881 BV=20 IBV=2e-05 CJO=2.0213e-10
	+VJ=0.386524 M=0.463886 FC=0.5 TT=1e-09
	+KF=0 AF=1
.ENDS






