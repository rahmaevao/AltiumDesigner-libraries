.SUBCKT BC846BLT1G C B E
	
	* Connections
		Q1 C B E Qbc846blt1g

	*modeles
		.MODEL Qbc846blt1g npn
		+IS=6.21868e-15 BF=313.939 NF=0.978615 VAF=808.652
		+IKF=0.0670247 ISE=6.72945e-10 NE=4 BR=31.3939
		+NR=1.03954 VAR=311.824 IKR=0.670247 ISC=5.02001e-14
		+NC=1.10677 RB=45.553 IRB=0.1 RBM=0.1
		+RE=0.18181 RC=0.909048 XTB=1.26632 XTI=1.16217
		+EG=1.206 CJE=7.31938e-12 VJE=0.479294 MJE=0.236218
		+TF=6.54085e-10 XTF=1000 VTF=8791.04 ITF=12.3428
		+CJC=1.97395e-12 VJC=0.95 MJC=0.33914 XCJC=1
		+FC=0.8 CJS=0 VJS=0.75 MJS=0.5
		+TR=1e-07 PTF=0 KF=0 AF=1

.ENDS BC846BLT1G
